class fifo_sb extends uvm_scoreboard;
`uvm_component_utils(fifo_sb)

function new(string name, uvm_component parent);
   super.new(name,parent);
endfunction
endclass
