/*********************************************************************************************************************************
 * Name                 : defines.sv
 * Creation Date        : 15-04-2022
 * Last Modified        : 09-05-2022
----------------------------------------------------------------------------------------------------------------------------------
 * Author               : Badam Mayur Krishna
 * Author's Email       : mayurkrishna.b@alpha-numero.tech
----------------------------------------------------------------------------------------------------------------------------------
* Description          :  Defines file for async_fifo project 
**********************************************************************************************************************************/

`define WIDTH 8
`define DEPTH 16

`define WRCLK_PERIOD 10
`define RDCLK_PERIOD 10


