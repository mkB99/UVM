
package fifo_pkg;

   import uvm_pkg::*;
   `include "uvm_macros.svh"

  `include "defines.sv"
  `include "wtrans.sv"
  `include "agent_config.sv"
  `include "wdrv.sv"
  `include "wmon.sv"
  `include "wseqr.sv"
  `include "wagent.sv"
  `include "wseqs.sv"
  `include "rtrans.sv"
  `include "rdrv.sv"
  `include "rmon.sv"
  `include "rseqr.sv"
  `include "rseqs.sv"
  `include "ragent.sv"
  `include "sb.sv"
  `include "env.sv"
  `include "fifo_base_test.sv"
  
endpackage
